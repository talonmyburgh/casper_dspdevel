-- megafunction wizard: %ROM: 1-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: ip_stratixiv_rom_r.vhd
-- Megafunction Name(s):
--      altsyncram
--
-- Simulation Library Files(s):
--      altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.0 Build 235 06/17/2009 SP 2 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2009 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY ip_stratixiv_rom_r IS
  GENERIC (
    g_adr_w     : NATURAL := 5;
    g_dat_w     : NATURAL := 8;
    g_nof_words : NATURAL := 2**5;
    g_init_file : STRING  := "UNUSED"
  );
  PORT (
    address   : IN STD_LOGIC_VECTOR(g_adr_w-1 DOWNTO 0);
    clock     : IN STD_LOGIC  := '1';
    clken     : IN STD_LOGIC  := '1';
    q         : OUT STD_LOGIC_VECTOR(g_dat_w-1 DOWNTO 0)
  );
END ip_stratixiv_rom_r;


ARCHITECTURE SYN OF ip_stratixiv_rom_r IS

  SIGNAL sub_wire0  : STD_LOGIC_VECTOR (g_dat_w-1 DOWNTO 0);

  COMPONENT altsyncram
  GENERIC (
    address_aclr_a    : STRING;
    clock_enable_input_a    : STRING;
    clock_enable_output_a   : STRING;
    init_file   : STRING;
    intended_device_family    : STRING;
    lpm_hint    : STRING;
    lpm_type    : STRING;
    numwords_a    : NATURAL;
    operation_mode    : STRING;
    outdata_aclr_a    : STRING;
    outdata_reg_a   : STRING;
    widthad_a   : NATURAL;
    width_a   : NATURAL;
    width_byteena_a   : NATURAL
  );
  PORT (
      clocken0  : IN STD_LOGIC ;
      clock0  : IN STD_LOGIC ;
      address_a : IN STD_LOGIC_VECTOR (g_adr_w-1 DOWNTO 0);
      q_a : OUT STD_LOGIC_VECTOR (g_dat_w-1 DOWNTO 0)
  );
  END COMPONENT;

BEGIN
  q    <= sub_wire0(g_dat_w-1 DOWNTO 0);

  altsyncram_component : altsyncram
  GENERIC MAP (
    address_aclr_a => "NONE",
    clock_enable_input_a => "NORMAL",
    clock_enable_output_a => "NORMAL",
    init_file => g_init_file,
    intended_device_family => "Stratix IV",
    lpm_hint => "ENABLE_RUNTIME_MOD=NO",
    lpm_type => "altsyncram",
    numwords_a => g_nof_words,
    operation_mode => "ROM",
    outdata_aclr_a => "NONE",
    outdata_reg_a => "CLOCK0",
    widthad_a => g_adr_w,
    width_a => g_dat_w,
    width_byteena_a => 1
  )
  PORT MAP (
    clocken0 => clken,
    clock0 => clock,
    address_a => address,
    q_a => sub_wire0
  );



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
-- Retrieval info: PRIVATE: AclrAddr NUMERIC "0"
-- Retrieval info: PRIVATE: AclrByte NUMERIC "0"
-- Retrieval info: PRIVATE: AclrOutput NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_ENABLE NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "9"
-- Retrieval info: PRIVATE: BlankMemory NUMERIC "0"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_A NUMERIC "1"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_A NUMERIC "1"
-- Retrieval info: PRIVATE: Clken NUMERIC "1"
-- Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
-- Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_A"
-- Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
-- Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
-- Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
-- Retrieval info: PRIVATE: MIFfilename STRING "fft_2n1024cos.hex"
-- Retrieval info: PRIVATE: NUMWORDS_A NUMERIC "32"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
-- Retrieval info: PRIVATE: RegAddr NUMERIC "1"
-- Retrieval info: PRIVATE: RegOutput NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: SingleClock NUMERIC "1"
-- Retrieval info: PRIVATE: UseDQRAM NUMERIC "0"
-- Retrieval info: PRIVATE: WidthAddr NUMERIC "5"
-- Retrieval info: PRIVATE: WidthData NUMERIC "18"
-- Retrieval info: PRIVATE: rden NUMERIC "0"
-- Retrieval info: CONSTANT: ADDRESS_ACLR_A STRING "NONE"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_A STRING "NORMAL"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_A STRING "NORMAL"
-- Retrieval info: CONSTANT: INIT_FILE STRING "fft_2n1024cos.hex"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: CONSTANT: LPM_HINT STRING "ENABLE_RUNTIME_MOD=NO"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
-- Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "32"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "ROM"
-- Retrieval info: CONSTANT: OUTDATA_ACLR_A STRING "NONE"
-- Retrieval info: CONSTANT: OUTDATA_REG_A STRING "CLOCK0"
-- Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "5"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "18"
-- Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
-- Retrieval info: USED_PORT: address 0 0 5 0 INPUT NODEFVAL address[4..0]
-- Retrieval info: USED_PORT: clken 0 0 0 0 INPUT VCC clken
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT VCC clock
-- Retrieval info: USED_PORT: q 0 0 18 0 OUTPUT NODEFVAL q[17..0]
-- Retrieval info: CONNECT: @address_a 0 0 5 0 address 0 0 5 0
-- Retrieval info: CONNECT: q 0 0 18 0 @q_a 0 0 18 0
-- Retrieval info: CONNECT: @clock0 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @clocken0 0 0 0 0 clken 0 0 0 0
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL ip_stratixiv_rom_r.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ip_stratixiv_rom_r.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ip_stratixiv_rom_r.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ip_stratixiv_rom_r.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ip_stratixiv_rom_r_inst.vhd FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ip_stratixiv_rom_r_waveforms.html TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL ip_stratixiv_rom_r_wave*.jpg FALSE
-- Retrieval info: LIB_FILE: altera_mf

--------------------------------------------------------------------------------
--
-- Copyright (C) 2016
-- ASTRON (Netherlands Institute for Radio Astronomy) <http://www.astron.nl/>
-- P.O.Box 2, 7990 AA Dwingeloo, The Netherlands
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
--------------------------------------------------------------------------------

-- Purpose: Multi-testbench for fil_ppf_wide using file data
-- Description:
--   Verify fil_ppf_wide using coefficients and data generated by
--   Matlab $RADIOHDL_WORK/applications/apertif/matlab/run_pfir.m
--   
-- Usage:
--   > as 4
--   > run -all

LIBRARY IEEE, common_pkg_lib;
USE IEEE.std_logic_1164.ALL;
USE common_pkg_lib.common_pkg.all;
USE work.fil_pkg.all;

ENTITY tb_tb_fil_ppf_wide_file_data IS
END tb_tb_fil_ppf_wide_file_data;

ARCHITECTURE tb OF tb_tb_fil_ppf_wide_file_data IS
  
  CONSTANT c_pipeline     : t_fil_ppf_pipeline := (1, 1, 1, 1, 1, 1, 0);
  
  CONSTANT c_coeff_prefix : string  := "hex/run_pfir_m_pfir_coeff_fircls1";
  CONSTANT c_data         : string  := "data/run_pfir_m_sinusoid_chirp_8b_16taps_128points_16b_16b.dat";  -- coefs, input and output data for 1 stream
  CONSTANT c_data15       : string  := "data/run_pfir_m_sinusoid_chirp_8b_15taps_128points_16b_16b.dat";  -- coefs, input and output data for 1 stream
 
  SIGNAL tb_end : STD_LOGIC := '0';  -- declare tb_end to avoid 'No objects found' error on 'when -label tb_end'
  
BEGIN

--g_big_endian_wb_in  : boolean := true;
--g_big_endian_wb_out : boolean := true;
--g_fil_ppf_pipeline : t_fil_ppf_pipeline := (1, 1, 1, 1, 1, 1, 0);
--  -- type t_fil_pipeline is record
--  --   -- generic for the taps and coefficients memory
--  --   mem_delay      : natural;  -- = 2
--  --   -- generics for the multiplier in in the filter unit
--  --   mult_input     : natural;  -- = 1
--  --   mult_product   : natural;  -- = 1
--  --   mult_output    : natural;  -- = 1
--  --   -- generics for the adder tree in in the filter unit
--  --   adder_stage    : natural;  -- = 1
--  --   -- generics for the requantizer in the filter unit
--  --   requant_remove_lsb : natural;  -- = 1
--  --   requant_remove_msb : natural;  -- = 0
--  -- end record;
--g_fil_ppf : t_fil_ppf := (1, 1, 64, 8, 1, 8, 20, 16);
--  -- type t_fil_ppf is record
--  --   wb_factor      : natural; -- = 1, the wideband factor
--  --   nof_chan       : natural; -- = default 0, defines the number of channels (=time-multiplexed input signals): nof channels = 2**nof_chan
--  --   nof_bands      : natural; -- = 128, the number of polyphase channels (= number of points of the FFT)
--  --   nof_taps       : natural; -- = 16, the number of FIR taps per subband
--  --   nof_streams    : natural; -- = 1, the number of streams that are served by the same coefficients.
--  --   backoff_w      : natural; -- = 0, number of bits for input backoff to avoid output overflow
--  --   in_dat_w       : natural; -- = 8, number of input bits per stream
--  --   out_dat_w      : natural; -- = 23, number of output bits (per stream). It is set to in_dat_w+coef_dat_w-1 = 23 to be sure the requantizer
--  --                                  does not remove any of the data in order to be able to verify with the original coefficients values.
--  --   coef_dat_w     : natural; -- = 16, data width of the FIR coefficients
--  -- end record;
--g_coefs_file_prefix   : string := "hex/run_pfir_m_pfir_coeff_fircls1";
--g_data_file           : string := "data/run_pfir_m_sinusoid_chirp_8b_16taps_128points_16b_16b.dat";  -- coefs, input and output data for 1 stream
--g_data_file_nof_lines : natural := 25600;  -- number of lines with input data that is available in the g_data_file
--g_data_file_nof_read  : natural := 5000;   -- number of lines with input data to read and simulate, must be <= g_data_file_nof_lines
--g_enable_in_val_gaps  : boolean := FALSE

  -- verify fil_ppf_wide for wb_factor=1, so effectively same as using fil_ppf_single directly
  u1_act                  : ENTITY work.tb_fil_ppf_wide_file_data GENERIC MAP (FALSE, FALSE, c_pipeline, (1, 0, 128, 16, 1, 1, 8, 16, 16), c_coeff_prefix, c_data,   25600, 25600, FALSE);
  u1_act_15taps           : ENTITY work.tb_fil_ppf_wide_file_data GENERIC MAP (FALSE, FALSE, c_pipeline, (1, 0, 128, 15, 1, 1, 8, 16, 16), c_coeff_prefix, c_data15, 25600,  5000, FALSE);
  u1_rnd                  : ENTITY work.tb_fil_ppf_wide_file_data GENERIC MAP (FALSE, FALSE, c_pipeline, (1, 0, 128, 16, 1, 1, 8, 16, 16), c_coeff_prefix, c_data,   25600,  5000, TRUE);
  u1_rnd_channels_streams : ENTITY work.tb_fil_ppf_wide_file_data GENERIC MAP (FALSE, FALSE, c_pipeline, (1, 1, 128, 16, 2, 1, 8, 16, 16), c_coeff_prefix, c_data,   25600,  5000, TRUE);
  
  -- verify fil_ppf_wide for wb_factor>1 (be = big endian, le = little endian)
  u4_act                  : ENTITY work.tb_fil_ppf_wide_file_data GENERIC MAP ( TRUE,  TRUE, c_pipeline, (4, 0, 128, 16, 1, 1, 8, 16, 16), c_coeff_prefix, c_data,   25600, 25600, FALSE);
  u4_act_be_le            : ENTITY work.tb_fil_ppf_wide_file_data GENERIC MAP ( TRUE, FALSE, c_pipeline, (4, 0, 128, 16, 1, 1, 8, 16, 16), c_coeff_prefix, c_data,   25600, 25600, FALSE);
  u4_act_le_be            : ENTITY work.tb_fil_ppf_wide_file_data GENERIC MAP (FALSE,  TRUE, c_pipeline, (4, 0, 128, 16, 1, 1, 8, 16, 16), c_coeff_prefix, c_data,   25600, 25600, FALSE);
  u4_act_le_le            : ENTITY work.tb_fil_ppf_wide_file_data GENERIC MAP (FALSE, FALSE, c_pipeline, (4, 0, 128, 16, 1, 1, 8, 16, 16), c_coeff_prefix, c_data,   25600, 25600, FALSE);
  u4_act_15taps           : ENTITY work.tb_fil_ppf_wide_file_data GENERIC MAP ( TRUE,  TRUE, c_pipeline, (4, 0, 128, 15, 1, 1, 8, 16, 16), c_coeff_prefix, c_data15, 25600,  5000, FALSE);
  u4_rnd                  : ENTITY work.tb_fil_ppf_wide_file_data GENERIC MAP ( TRUE,  TRUE, c_pipeline, (4, 0, 128, 16, 1, 1, 8, 16, 16), c_coeff_prefix, c_data,   25600,  5000, TRUE);
  u4_rnd_channels_streams : ENTITY work.tb_fil_ppf_wide_file_data GENERIC MAP ( TRUE,  TRUE, c_pipeline, (4, 1, 128, 16, 4, 1, 8, 16, 16), c_coeff_prefix, c_data,   25600,  5000, TRUE);

END tb;

-------------------------------------------------------------------------------
--
-- Copyright 2020
-- ASTRON (Netherlands Institute for Radio Astronomy) <http://www.astron.nl/>
-- P.O.Box 2, 7990 AA Dwingeloo, The Netherlands
-- 
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
-- 
--     http://www.apache.org/licenses/LICENSE-2.0
-- 
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-------------------------------------------------------------------------------

LIBRARY IEEE, common_pkg_lib, common_components_lib, technology_lib;
USE IEEE.std_logic_1164.ALL;
USE common_pkg_lib.common_pkg.ALL;
USE work.tech_mult_component_pkg.all;
USE technology_lib.technology_select_pkg.ALL;

ENTITY tech_complex_mult IS
	GENERIC(
		g_sim              : BOOLEAN := TRUE;
		g_sim_level        : NATURAL := 0; -- 0: Simulate variant passed via g_use_variant for given technology
		g_use_variant      : STRING  := "4DSP";
		g_use_dsp          : STRING  := "YES"; --! Implement multiplications in DSP48 or not
		g_in_a_w           : POSITIVE;
		g_in_b_w           : POSITIVE;
		g_out_p_w          : POSITIVE;  -- default use g_out_p_w = g_in_a_w+g_in_b_w = c_prod_w
		g_conjugate_b      : BOOLEAN := FALSE;
		g_pipeline_input   : NATURAL := 1; -- 0 or 1
		g_pipeline_product : NATURAL := 0; -- 0 or 1
		g_pipeline_adder   : NATURAL := 1; -- 0 or 1
		g_pipeline_output  : NATURAL := 1 -- >= 0
	);
	PORT(
		rst       : IN  STD_LOGIC := '0';
		clk       : IN  STD_LOGIC;
		clken     : IN  STD_LOGIC := '1';
		in_ar     : IN  STD_LOGIC_VECTOR(g_in_a_w - 1 DOWNTO 0);
		in_ai     : IN  STD_LOGIC_VECTOR(g_in_a_w - 1 DOWNTO 0);
		in_br     : IN  STD_LOGIC_VECTOR(g_in_b_w - 1 DOWNTO 0);
		in_bi     : IN  STD_LOGIC_VECTOR(g_in_b_w - 1 DOWNTO 0);
		result_re : OUT STD_LOGIC_VECTOR(g_out_p_w - 1 DOWNTO 0);
		result_im : OUT STD_LOGIC_VECTOR(g_out_p_w - 1 DOWNTO 0)
	);
END tech_complex_mult;

ARCHITECTURE str of tech_complex_mult is

	--! Force to maximum 18 bit width, because:
	--! . the ip_cmult_infer is generated for 18b inputs and 36b output and then uses 4 real multipliers and no additional registers
	--! . if one input   > 18b then another IP needs to be regenerated and that will use  8 real multipliers and some extra LUTs and registers
	--! . if both inputs > 18b then another IP needs to be regenerated and that will use 16 real multipliers and some extra LUTs and registers
	--! . if the output is set to 18b+18b + 1b =37b to account for the sum then another IP needs to be regenerated and that will use some extra registers
	--! ==> for inputs <= 18b this ip_complex_mult is appropriate and it can not be made parametrisable to fit also inputs > 18b.

	-- sim_model=1
	SIGNAL result_re_undelayed : STD_LOGIC_VECTOR(g_in_b_w + g_in_a_w - 1 DOWNTO 0);
	SIGNAL result_im_undelayed : STD_LOGIC_VECTOR(g_in_b_w + g_in_a_w - 1 DOWNTO 0);

begin

	gen_ip_xpm_rtl_4dsp : IF c_tech_select_default = c_tech_xpm AND g_use_variant = "4DSP" GENERATE  -- Xilinx
		u1 : ip_cmult_rtl_4dsp
			generic map(
				g_use_dsp          => g_use_dsp,
				g_in_a_w           => g_in_a_w,
				g_in_b_w           => g_in_b_w,
				g_out_p_w          => g_out_p_w,
				g_conjugate_b      => g_conjugate_b,
				g_pipeline_input   => g_pipeline_input,
				g_pipeline_product => g_pipeline_product,
				g_pipeline_adder   => g_pipeline_adder,
				g_pipeline_output  => g_pipeline_output
			)
			port map(
				rst       => rst,
				clk       => clk,
				clken     => clken,
				in_ar     => in_ar,
				in_ai     => in_ai,
				in_br     => in_br,
				in_bi     => in_bi,
				result_re => result_re,
				result_im => result_im
			);
	end generate;

	gen_ip_xpm_rtl_3dsp : IF c_tech_select_default = c_tech_xpm AND g_use_variant = "3DSP" GENERATE  -- Xilinx
		u1 : ip_cmult_rtl_3dsp
			generic map(
				g_use_dsp          => g_use_dsp,
				g_in_a_w           => g_in_a_w,
				g_in_b_w           => g_in_b_w,
				g_out_p_w          => g_out_p_w,
				g_conjugate_b      => g_conjugate_b,
				g_pipeline_input   => g_pipeline_input,
				g_pipeline_product => g_pipeline_product,
				g_pipeline_adder   => g_pipeline_adder,
				g_pipeline_output  => g_pipeline_output
			)
			port map(
				rst       => rst,
				clk       => clk,
				clken     => clken,
				in_ar     => in_ar,
				in_ai     => in_ai,
				in_br     => in_br,
				in_bi     => in_bi,
				result_re => result_re,
				result_im => result_im
			);
	end generate;

	-------------------------------------------------------------------------------
	-- Model: forward concatenated inputs to the 'result' output
	-- 
	-- Example:
	--                                    ______ 
	-- Input B.real (in_br) = 0x1111 --> |      |
	--        .imag (in_bi) = 0xBBBB --> |      |
	--                                   | mult | --> Output result.real = 0x11110000
	-- Input A.real (in_ar) = 0x0000 --> |      |                  .imag = 0xBBBBAAAA
	--        .imag (in_ai) = 0xAAAA --> |______|
	-- 
	-- Note: this model is synthsizable as well.
	-- 
	-------------------------------------------------------------------------------
	gen_sim_level_1 : IF g_sim = TRUE AND g_sim_level = 1 GENERATE --FIXME: g_sim required? This is synthesizable.

		result_re_undelayed <= in_br & in_ar;
		result_im_undelayed <= in_bi & in_ai;

		u_common_pipeline_re : entity common_components_lib.common_pipeline
			generic map(
				g_pipeline  => 3,
				g_in_dat_w  => g_in_b_w + g_in_a_w,
				g_out_dat_w => g_out_p_w
			)
			port map(
				clk     => clk,
				in_dat  => result_re_undelayed,
				out_dat => result_re
			);

		u_common_pipeline_im : entity common_components_lib.common_pipeline
			generic map(
				g_pipeline  => 3,
				g_in_dat_w  => g_in_b_w + g_in_a_w,
				g_out_dat_w => g_out_p_w
			)
			port map(
				clk     => clk,
				in_dat  => result_im_undelayed,
				out_dat => result_im
			);

	END GENERATE;
end str;

-- author: Auguust 2023 - Andrew Martens but compiled from Astron sources with improvements mostly to reduce BRAM use 
-- add sync functionality and improve timing

library IEEE, common_pkg_lib, casper_ram_lib, casper_multiplier_lib, casper_adder_lib, casper_requantize_lib, technology_lib;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;
use common_pkg_lib.common_pkg.ALL;
use casper_ram_lib.common_ram_pkg.ALL;
use technology_lib.technology_select_pkg.ALL;
use work.pfb_fir_pkg.ALL;

entity pfb_fir is
  generic (
    g_coefs_file    : string             := c_pfb_fir_coefs_file; --! coefficients file generated by fil_ppf_create.py
    g_ram_primitive : string             := "auto";
    g_pfb_fir       : t_pfb_fir          := c_pfb_fir          		-- standard record from package
  );
  port (
    clk       : in std_logic;    
    sync_in   : in std_logic;
    din       : in t_pfb_fir_array_in((g_pfb_fir.wb_factor*g_pfb_fir.n_streams)-1 downto 0);
    en        : in std_logic;
    sync_out  : out std_logic;
    dout      : out t_pfb_fir_array_out((g_pfb_fir.wb_factor*g_pfb_fir.n_streams)-1 downto 0);
    dvalid    : out std_logic
  );
end pfb_fir;

architecture rtl of pfb_fir is
-- control logic

  constant c_tap_length         : natural := (g_pfb_fir.n_bins/g_pfb_fir.wb_factor)*(2**g_pfb_fir.n_chans);
  constant c_addr_w             : natural := ceil_log2(c_tap_length);
  signal master_counter         : std_logic_vector(c_addr_w-1 downto 0);
  
  -- note that this differs from Astron's delay. 
  constant c_sync_delay         : natural := c_tap_length * (g_pfb_fir.n_taps-1); 
  signal sync_cnt               : std_logic_vector(ceil_log2(c_sync_delay)-1 downto 0);
  signal sync_out_int           : std_logic;
  signal dvalid_int             : std_logic;
  signal dout_int               : t_pfb_fir_array_out((g_pfb_fir.wb_factor*g_pfb_fir.n_streams)-1 downto 0);
  
  constant c_delay_adder_tree   : natural := ceil_log2(g_pfb_fir.n_taps) * g_pfb_fir.add_latency;
  constant c_delay_total        : natural := g_pfb_fir.mem_latency + g_pfb_fir.mult_latency + c_delay_adder_tree + g_pfb_fir.conv_latency;
      
  signal en_delay               : std_logic_vector(c_delay_total-1 downto 0) := (others => '0');           -- enable pipeline
  signal sync_in_delay          : std_logic_vector(c_delay_total-1 downto 0) := (others => '0');
  
-- coefficients
  constant c_coefs_total                : natural   := g_pfb_fir.wb_factor * g_pfb_fir.n_taps;
  constant c_coef_mem_addr_w            : natural   := c_addr_w - g_pfb_fir.n_chans;
  constant c_coef_mem_data_w            : natural   := g_pfb_fir.coef_w;
  constant c_coefs_postfix              : string    := sel_a_b(c_tech_select_default = c_tech_xpm, ".mem", ".mif");                                                                                                    
  constant c_coef_mem                   : t_c_mem   := (latency   => g_pfb_fir.mem_latency,
                                              adr_w     => c_coef_mem_addr_w,
                                              dat_w     => c_coef_mem_data_w,
                                              nof_dat   => g_pfb_fir.n_bins,
                                              init_sl   => '0');  -- use '0' instead of 'X' to avoid RTL RAM simulation warnings due to read before write
  signal coef_rdaddr, coef_rdaddr_inv   : std_logic_vector(c_coef_mem_addr_w-1 downto 0);     
  TYPE t_coef_array is array (integer range <>) of std_logic_vector(c_coef_mem_data_w-1 DOWNTO 0);
  signal coef_vec                       : t_coef_array(c_coefs_total-1 downto 0) := (others => (others => '0'));
  
-- taps 
  constant c_tap_data_w                 : natural := g_pfb_fir.wb_factor * g_pfb_fir.n_streams * g_pfb_fir.din_w;
  constant c_taps_mem_data_w            : natural := c_tap_data_w * (g_pfb_fir.n_taps-1);
  constant c_taps_mem                   : t_c_mem   := (latency   => g_pfb_fir.mem_latency,
                                              adr_w     => c_addr_w,
                                              dat_w     => c_taps_mem_data_w,
                                              nof_dat   => (g_pfb_fir.n_bins/g_pfb_fir.wb_factor)*(2**g_pfb_fir.n_chans),
                                              init_sl   => '0');  -- use '0' instead of 'X' to avoid RTL RAM simulation warnings due to read before write
  signal taps_wren                      : std_logic := '0';
  type   t_in_dat_delay is array (g_pfb_fir.mem_latency-1 downto 0) of std_logic_vector(c_tap_data_w-1 downto 0);
  signal din_delay                      : t_in_dat_delay;
  
  signal taps_rdaddr, taps_wraddr       : std_logic_vector(c_addr_w-1 downto 0);
  signal taps_in_vec, taps_out_vec      : std_logic_vector(c_taps_mem_data_w-1 downto 0) := (others => '0'); 
  
      
--multipliers
  constant c_mult_din_w     : natural := g_pfb_fir.padding + g_pfb_fir.din_w;        -- add optional input padding to fit output overshoot
  constant c_prod_w         : natural := g_pfb_fir.din_w + g_pfb_fir.coef_w - 1;    -- skip double sign bit
  constant c_n_mults        : natural := g_pfb_fir.wb_factor * g_pfb_fir.n_taps * g_pfb_fir.n_streams;

  signal mult_din, mult_din_reordered : std_logic_vector(c_n_mults * g_pfb_fir.din_w-1 downto 0); 
  signal mult_din_padding             : std_logic_vector(c_n_mults * c_mult_din_w-1 downto 0);  -- taps input data with padding 
  signal prod_vec                     : std_logic_vector(c_n_mults * c_prod_w-1 downto 0);
                                              
--adder tree  
  constant c_gain_w         : natural := 0;   -- no need for adder bit growth so fixed 0, because filter coefficients should have DC gain <= 1.
                                              -- The adder tree bit growth depends on DC gain of FIR coefficients, not on ceil_log2(g_fil_ppf.nof_taps). 
  constant c_sum_w          : natural := c_prod_w + c_gain_w;
  constant c_ppf_lsb_w      : natural := c_sum_w - g_pfb_fir.dout_w;
  
  signal adder_out          : std_logic_vector(g_pfb_fir.wb_factor*c_sum_w-1 downto 0) := (others => '0');
  
--requantisation  
  signal requant_out        : std_logic_vector(g_pfb_fir.wb_factor*g_pfb_fir.dout_w-1 downto 0); 
       
begin

-- control of addresses, pipelines etc
proc_master: process(clk) begin 
  if rising_edge(clk) then --everything is synchronous 
    if (sync_in = '1') then
      master_counter <= (others => '0');
    else 
      if (en = '1') then
        master_counter <= std_logic_vector(unsigned(master_counter) + 1);
      end if;
    end if; 
    
    -- enable pipeline
    en_delay(0) <= en;
    en_delay(c_delay_total-1 downto 1) <= en_delay(c_delay_total-2 downto 0);  
    
    --sync pipeline
    sync_in_delay(0) <= sync_in;
    sync_in_delay(c_delay_total-1 downto 1) <= sync_in_delay(c_delay_total-2 downto 0);

    --sync counter
    if (sync_in_delay(c_delay_total-1) = '1') then
      sync_cnt <= (others => '0');
    else 
      -- increment the sync counter if counting and a value is passing
      if (unsigned(sync_cnt) < c_sync_delay and en_delay(c_delay_total-1) = '1') then
        sync_cnt <= std_logic_vector(unsigned(sync_cnt) + 1);
      end if;
    end if;
    
    --generate a sync out on the last value
    if(unsigned(sync_cnt) = (c_sync_delay-1) and en_delay(c_delay_total-1) = '1') then
      sync_out_int <= '1';
    else 
      sync_out_int <= '0';
    end if;
    
    dvalid_int <= en_delay(c_delay_total-1);
    
  end if; --rising_edge(clk)
end process proc_master;

dvalid <= dvalid_int;
sync_out <= sync_out_int;
dout <= dout_int;

-- taps
proc_taps:process(clk) begin
  if(rising_edge(clk)) then
    din_delay(0) <= din(0); 
    din_delay(g_pfb_fir.mem_latency-1 downto 1) <= din_delay(g_pfb_fir.mem_latency-2 downto 0);
   
    -- the write address is delayed while we wait for the data from the read 
    if(sync_in_delay(g_pfb_fir.mem_latency-1) = '1') then
      taps_wraddr <= (others => '0');
    else
      if(en_delay(g_pfb_fir.mem_latency-1) = '1') then
        taps_wraddr <= std_logic_vector(unsigned(taps_wraddr) + 1);
      end if;
    end if;
  end if;
end process;    

taps_rdaddr <= master_counter(c_addr_w-1 downto 0); --lsbs for channels too
-- we feed new data in from the least significant bits
taps_in_vec(c_taps_mem_data_w-1 downto 0) <=  taps_out_vec(c_taps_mem_data_w-c_tap_data_w-1 downto 0) & din_delay(g_pfb_fir.mem_latency-1);
taps_wren <= en_delay(g_pfb_fir.mem_latency-1);

u_taps_mem : entity casper_ram_lib.common_ram_r_w                                                          
  generic map (                                                                                    
    g_ram           => c_taps_mem,                                                                           
    g_init_file     => "UNUSED",     -- assume block RAM gets initialized to '0' by default in simulation
    g_ram_primitive => g_ram_primitive
  )                                                                                               
  port map (                                                                                                                                                                     
    clk       => clk,
    clken     => '1',                                                                               
    wr_en     => taps_wren,                                                                              
    wr_adr    => taps_wraddr,                                                                            
    wr_dat    => taps_in_vec,                                                                            
    rd_en     => '1',                                                                               
    rd_adr    => taps_rdaddr,                                                                            
    rd_dat    => taps_out_vec,  
    rd_val    => open                                                                               
  );  

-- coefficients

coef_rdaddr <= master_counter(c_addr_w-1 downto g_pfb_fir.n_chans);
coef_rdaddr_inv <= not(coef_rdaddr);

gen_coefs: for I in 0 to g_pfb_fir.wb_factor-1 generate
begin
  gen_coeffs: for C in 0 to (g_pfb_fir.n_taps/2)-1 generate
    constant c_coef_offset        : natural := I * g_pfb_fir.n_taps/2 + C; --base offset in output vector
  begin
    u_coef_mem : entity casper_ram_lib.common_rom_r_r
      generic map (
        g_ram           =>     c_coef_mem,
        g_init_file     =>     sel_a_b(g_coefs_file = "UNUSED", 
                               g_coefs_file, 
                               g_coefs_file 
                               & "_" & integer'image(g_pfb_fir.wb_factor) 
                               & "wb" & "_" 
                               & NATURAL'IMAGE((I * g_pfb_fir.n_taps) + C) & c_coefs_postfix),
        g_ram_primitive =>     g_ram_primitive,
        g_true_dual_port =>    TRUE
      ) 
      port map 
      (
        clk =>        clk,
        clken =>      '1',
        adr_a =>      coef_rdaddr, 
        rd_en_a =>    '1',
        rd_dat_a =>   coef_vec(c_coef_offset),
        rd_val_a =>   open,
        adr_b =>      coef_rdaddr_inv, --count backwards on other port
        rd_en_b =>    '1',
        rd_dat_b =>   coef_vec(c_coefs_total-c_coef_offset-1) --coefficients are symmetrical
      );
  end generate; -- Coeffs
end generate; --I     

--multipliers 
 
--we get the tap with delay 0 for (almost) free
mult_din((c_n_mults * g_pfb_fir.din_w)-1 downto 0) <= taps_out_vec & din_delay(g_pfb_fir.mem_latency-1);
  
gen_mults: for I in 0 to g_pfb_fir.wb_factor-1 generate
begin
  gen_taps: for T in 0 to g_pfb_fir.n_taps-1 generate
    constant c_coef_offset : natural := (I * g_pfb_fir.n_taps) + T;
  begin
    gen_streams: for S in 0 to g_pfb_fir.n_streams-1 generate
      constant c_src_offset: natural := T * (g_pfb_fir.wb_factor * g_pfb_fir.n_streams) + (I * g_pfb_fir.n_streams) + S;
      constant c_dest_offset : natural := (I * g_pfb_fir.n_streams * g_pfb_fir.n_taps) + (S * g_pfb_fir.n_taps) + T;  
    begin       
      mult_din_reordered(((c_dest_offset+1)*g_pfb_fir.din_w)-1 downto c_dest_offset*g_pfb_fir.din_w) <= mult_din(((c_src_offset+1)*g_pfb_fir.din_w)-1 downto c_src_offset*g_pfb_fir.din_w);

      mult_din_padding((c_dest_offset+1)*c_mult_din_w-1 downto c_dest_offset*c_mult_din_w) <= resize_svec(mult_din((c_dest_offset+1)*g_pfb_fir.din_w-1 downto c_dest_offset*g_pfb_fir.din_w), c_mult_din_w);
    
      u_multiplier : entity casper_multiplier_lib.common_mult
      generic map (
        g_use_dsp          => "YES",
        g_in_a_w           => c_mult_din_w,   
        g_in_b_w           => g_pfb_fir.coef_w, 
        g_out_p_w          => c_prod_w,                              
        g_pipeline_input   => sel_a_b(g_pfb_fir.mult_latency > 2, 1, 0),
        g_pipeline_product => sel_a_b(g_pfb_fir.mult_latency > 2, 1, 0),  
        g_pipeline_output  => sel_a_b(g_pfb_fir.mult_latency > 2, g_pfb_fir.mult_latency-2, g_pfb_fir.mult_latency)       
      )
      port map (
        rst      => '0',
        clk      => clk,
        clken    => '1',
        in_a     => mult_din_padding((c_dest_offset+1)*c_mult_din_w-1 downto c_dest_offset*c_mult_din_w),
        in_b     => coef_vec(c_coef_offset),
        result   => prod_vec((c_dest_offset+1)*c_prod_w-1 downto c_dest_offset*c_prod_w)
      );
    
    end generate;
  end generate; -- T 
end generate; -- I  

--adder trees
gen_add_quantise: for I in 0 to g_pfb_fir.wb_factor-1 generate
begin
    gen_streams: for S in 0 to g_pfb_fir.n_streams-1 generate
      constant c_offset : natural := (I * g_pfb_fir.n_streams) + S;
    begin
    
      u_adder_tree : entity casper_adder_lib.common_adder_tree 
      generic map (
        g_representation => "SIGNED",
        g_pipeline       => g_pfb_fir.add_latency,          
        g_nof_inputs     => g_pfb_fir.n_taps,
        g_dat_w          => c_prod_w,
        g_sum_w          => c_sum_w 
      )
      port map (
        clk    => clk,
        in_dat => prod_vec((c_offset+1)*g_pfb_fir.n_taps*c_prod_w-1 downto c_offset*g_pfb_fir.n_taps*c_prod_w),
        sum    => adder_out((c_offset+1)*c_sum_w-1 downto c_offset*c_sum_w)
      );

--requantisation
      
      u_requantize : entity casper_requantize_lib.common_requantize
      generic map (
        g_representation      => "SIGNED",      
        g_lsb_w               => c_ppf_lsb_w,  
        g_lsb_round           => TRUE,           
        g_lsb_round_clip      => FALSE,      
        g_msb_clip            => FALSE,            
        g_msb_clip_symmetric  => FALSE,  
        g_pipeline_remove_lsb => 1, --hardcoded for now 
        g_pipeline_remove_msb => 0, --hardcoded for now
        g_in_dat_w            => c_sum_w,            
        g_out_dat_w           => g_pfb_fir.dout_w
      )
      port map (
        clk        => clk,
        clken      => '1',
        in_dat     => adder_out(((c_offset+1)*c_sum_w)-1 downto c_offset*c_sum_w),
        out_dat    => requant_out(((c_offset+1)*g_pfb_fir.dout_w)-1 downto c_offset*g_pfb_fir.dout_w), 
        out_ovr    => open
      );         
      
      --register the outputs to align with sync and dvalid
      process(clk) begin
        if(rising_edge(clk)) then
          dout_int(c_offset) <= requant_out(((c_offset+1)*g_pfb_fir.dout_w)-1 downto c_offset*g_pfb_fir.dout_w);
        end if;
      end process;
                   
    end generate; --S 
end generate; --I

end rtl;
